library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity displaybuffer is
    generic (
        OBJECT_SIZE : natural := 16;
        PIXEL_SIZE : natural := 24;
        RES_X : natural := 1280;
        RES_Y : natural := 720
    );
    port (
		S_AXI_ACLK		   : in std_logic;
        video_active       : in  std_logic;
        pixel_x, pixel_y   : in  std_logic_vector(OBJECT_SIZE-1 downto 0);
        object1x, object1y : in  std_logic_vector(OBJECT_SIZE-1 downto 0);
        object2x, object2y : in  std_logic_vector(OBJECT_SIZE-1 downto 0);
        backgrnd_rgb       : in  std_logic_vector(PIXEL_SIZE-1 downto 0);
        rgb                : out std_logic_vector(PIXEL_SIZE-1 downto 0)
    );
end displaybuffer;

architecture rtl of displaybuffer is
    -- create a 5 pixel vertical wall
--    constant WALL_X_L: integer := 60;
--    constant WALL_X_R: integer := 65;

    -- 1st object is a vertical box 48x8 pixel
--    constant BOX_SIZE_X: integer :=  8;
--    constant BOX_SIZE_Y: integer := 48;
    -- x, y coordinates of the box
--    signal box_x_l : unsigned (OBJECT_SIZE-1 downto 0);
--    signal box_y_t : unsigned (OBJECT_SIZE-1 downto 0);
--    signal box_x_r : unsigned (OBJECT_SIZE-1 downto 0);
--    signal box_y_b : unsigned (OBJECT_SIZE-1 downto 0);

    -- 2nd object is a ball
    constant BALL_SIZE_8 : integer := 8;
    type rom_type_8 is array ( 0 to 7 ) of std_logic_vector( 7 downto 0 );
    constant BALL_ROM_8: rom_type_8 := (
       "00111100",
       "01111110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111110",
       "00111100"
    );
	
	constant BALL_SIZE_32 : integer := 32;
    type rom_type_32 is array ( 0 to 31 ) of std_logic_vector( 31 downto 0 );
    constant BALL_ROM_32: rom_type_32 := (
       "00000000000111111111100000000000",
       "00000000111111111111111100000000",
       "00000001111111111111111110000000",
       "00000111111111111111111111100000",
       "00001111111111111111111111110000",
       "00011111111111111111111111111000",
       "00011111111111111111111111111000",
       "00111111111111111111111111111100",
       "01111111111111111111111111111110",
       "01111111111111111111111111111110",
       "01111111111111111111111111111110",
       "11111111111111111111111111111111",
       "11111111111111111111111111111111",
       "11111111111111111111111111111111",
       "11111111111111111111111111111111",
       "11111111111111111111111111111111",
       "11111111111111111111111111111111",
       "11111111111111111111111111111111",
       "11111111111111111111111111111111",
       "11111111111111111111111111111111",
       "11111111111111111111111111111111",
       "01111111111111111111111111111110",
       "01111111111111111111111111111110",
       "01111111111111111111111111111110",
       "00111111111111111111111111111100",
       "00011111111111111111111111111000",
       "00011111111111111111111111111000",
       "00001111111111111111111111110000",
       "00000111111111111111111111100000",
       "00000001111111111111111110000000",
       "00000000111111111111111100000000",
       "00000000000111111111100000000000"
    );
	
	type BALL32_COLOR_TYPE is array ( 0 to BALL_SIZE_32 - 1, 0 to  BALL_SIZE_32 - 1 ) of integer;
	
	constant BALL32_COLOR : BALL32_COLOR_TYPE := (
		( 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 167, 172, 174, 177, 179, 181, 182, 183, 183, 183, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255, 255 ),
		( 255, 255, 255, 255, 255, 255, 255, 255, 174, 165, 169, 172, 176, 179, 182, 184, 186, 187, 188, 188, 188, 188, 187, 181, 255, 255, 255, 255, 255, 255, 255, 255 ),
		( 255, 255, 255, 255, 255, 255, 255, 162, 162, 168, 173, 178, 181, 185, 188, 191, 193, 194, 195, 195, 195, 194, 192, 190, 188, 255, 255, 255, 255, 255, 255, 255 ),
		( 255, 255, 255, 255, 255, 255, 150, 154, 161, 170, 178, 182, 186, 189, 193, 197, 199, 200, 202, 202, 201, 200, 198, 196, 193, 190, 177, 255, 255, 255, 255, 255 ),
		( 255, 255, 255, 255, 255, 137, 144, 153, 163, 172, 179, 186, 191, 195, 199, 202, 205, 206, 208, 208, 207, 206, 204, 202, 199, 194, 190, 184, 255, 255, 255, 255 ),
		( 255, 255, 255, 255, 122, 132, 143, 154, 164, 173, 181, 189, 195, 200, 204, 208, 210, 213, 214, 214, 214, 212, 209, 207, 204, 199, 194, 190, 184, 255, 255, 255 ),
		( 255, 255, 255, 111, 119, 131, 144, 155, 165, 174, 182, 191, 198, 203, 209, 213, 216, 219, 220, 220, 220, 218, 215, 212, 208, 204, 199, 193, 189, 255, 255, 255 ),
		( 255, 255, 102, 107, 118, 131, 143, 154, 165, 174, 184, 192, 199, 207, 213, 218, 222, 224, 226, 226, 226, 224, 221, 217, 213, 208, 202, 197, 191, 186, 255, 255 ),
		( 255, 255, 99, 103, 116, 129, 142, 153, 164, 175, 184, 193, 201, 209, 216, 222, 226, 230, 232, 233, 232, 229, 225, 221, 217, 211, 205, 200, 194, 188, 179, 255 ),
		( 255, 93, 95, 101, 114, 127, 140, 152, 163, 175, 184, 194, 203, 211, 218, 225, 230, 236, 238, 239, 238, 234, 230, 225, 219, 214, 208, 202, 196, 190, 184, 255 ),
		( 255, 88, 90, 99, 112, 124, 138, 150, 162, 174, 184, 194, 203, 212, 220, 227, 234, 240, 244, 245, 244, 239, 234, 228, 222, 216, 209, 204, 198, 191, 185, 174 ),
		( 81, 83, 86, 94, 108, 122, 135, 148, 160, 171, 182, 193, 202, 211, 220, 227, 235, 242, 249, 252, 248, 242, 236, 229, 223, 217, 211, 205, 198, 192, 185, 180 ),
		( 76, 78, 82, 90, 104, 118, 132, 144, 156, 168, 180, 191, 201, 210, 219, 227, 235, 242, 249, 253, 249, 242, 236, 229, 223, 217, 211, 205, 198, 192, 185, 180 ),
		( 72, 75, 79, 86, 99, 113, 127, 140, 152, 165, 177, 187, 198, 208, 216, 224, 232, 239, 244, 245, 244, 240, 234, 228, 222, 216, 209, 204, 198, 191, 184, 179 ),
		( 67, 71, 75, 82, 95, 107, 121, 135, 148, 160, 172, 183, 193, 203, 213, 220, 227, 234, 238, 239, 238, 235, 231, 226, 220, 214, 208, 202, 196, 190, 183, 178 ),
		( 63, 66, 70, 75, 88, 102, 115, 128, 143, 154, 166, 177, 187, 197, 206, 214, 221, 226, 230, 231, 231, 229, 226, 222, 217, 211, 205, 200, 195, 189, 182, 176 ),
		( 59, 62, 67, 70, 81, 95, 109, 122, 135, 147, 159, 171, 181, 191, 199, 207, 213, 219, 221, 223, 223, 222, 220, 217, 213, 208, 203, 198, 192, 186, 180, 175 ),
		( 55, 58, 63, 66, 74, 88, 101, 114, 127, 139, 150, 163, 173, 183, 191, 199, 205, 210, 213, 215, 216, 215, 213, 211, 208, 204, 199, 194, 189, 183, 177, 172 ),
		( 50, 54, 58, 63, 68, 79, 92, 106, 119, 131, 143, 153, 164, 174, 182, 189, 195, 200, 204, 206, 207, 207, 205, 204, 201, 198, 195, 190, 185, 180, 174, 169 ),
		( 46, 50, 55, 58, 62, 71, 84, 97, 109, 121, 133, 143, 153, 164, 172, 179, 185, 190, 194, 196, 197, 198, 197, 196, 194, 192, 190, 186, 182, 177, 171, 167 ),
		( 43, 46, 51, 54, 58, 64, 75, 88, 99, 111, 122, 134, 143, 153, 161, 168, 174, 180, 183, 186, 188, 189, 189, 188, 186, 184, 182, 181, 178, 173, 168, 163 ),
		( 38, 42, 46, 50, 54, 58, 65, 77, 88, 101, 111, 122, 132, 141, 149, 157, 163, 168, 172, 175, 177, 178, 179, 179, 178, 176, 175, 174, 171, 168, 164, 255 ),
		( 255, 38, 42, 46, 50, 54, 58, 66, 78, 90, 100, 110, 120, 129, 137, 144, 151, 156, 160, 164, 166, 168, 169, 169, 169, 168, 167, 166, 164, 163, 159, 255 ),
		( 255, 34, 37, 42, 47, 50, 54, 58, 67, 77, 88, 98, 107, 116, 124, 131, 138, 143, 148, 151, 154, 156, 157, 158, 159, 159, 158, 157, 156, 154, 146, 255 ),
		( 255, 0, 35, 38, 42, 46, 51, 54, 58, 66, 76, 86, 95, 103, 111, 118, 124, 130, 135, 138, 142, 145, 146, 147, 148, 148, 147, 147, 146, 144, 255, 255 ),
		( 255, 255, 30, 34, 38, 42, 46, 50, 54, 58, 63, 73, 82, 91, 98, 105, 111, 117, 122, 126, 129, 132, 134, 135, 136, 136, 136, 136, 136, 134, 255, 255 ),
		( 255, 255, 255, 31, 34, 38, 42, 46, 50, 54, 58, 62, 68, 77, 84, 91, 98, 103, 108, 113, 116, 119, 120, 123, 124, 124, 124, 126, 129, 255, 255, 255 ),
		( 255, 255, 255, 255, 30, 34, 38, 42, 46, 50, 54, 58, 62, 65, 72, 77, 83, 89, 93, 98, 102, 105, 107, 109, 111, 114, 117, 121, 255, 255, 255, 255 ),
		( 255, 255, 255, 255, 255, 31, 34, 38, 42, 46, 50, 54, 58, 61, 65, 70, 74, 78, 82, 86, 90, 94, 98, 102, 105, 110, 115, 255, 255, 255, 255, 255 ),
		( 255, 255, 255, 255, 255, 255, 30, 34, 37, 41, 46, 50, 54, 58, 62, 66, 70, 74, 78, 81, 85, 90, 93, 98, 103, 106, 255, 255, 255, 255, 255, 255 ),
		( 255, 255, 255, 255, 255, 255, 255, 26, 34, 38, 41, 45, 49, 54, 57, 61, 65, 69, 74, 77, 81, 85, 90, 95, 91, 255, 255, 255, 255, 255, 255, 255 ),
		( 255, 255, 255, 255, 255, 255, 255, 255, 255, 32, 39, 42, 46, 49, 54, 58, 62, 66, 70, 74, 78, 83, 84, 255, 255, 255, 255, 255, 255, 255, 255, 255 )
	);
	
	constant BALL32_ALPHA : BALL32_COLOR_TYPE := (
		( 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 26, 43, 59, 65, 69, 72, 61, 43, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ),
		( 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 30, 46, 57, 64, 71, 77, 82, 85, 87, 89, 85, 67, 36, 4, 0, 0, 0, 0, 0, 0, 0, 0 ),
		( 0, 0, 0, 0, 0, 0, 0, 6, 29, 42, 51, 61, 70, 79, 86, 93, 98, 102, 105, 105, 105, 106, 103, 83, 33, 0, 0, 0, 0, 0, 0, 0 ),
		( 0, 0, 0, 0, 0, 0, 14, 42, 52, 56, 63, 72, 82, 92, 100, 107, 113, 117, 120, 121, 120, 117, 112, 109, 104, 60, 2, 0, 0, 0, 0, 0 ),
		( 0, 0, 0, 0, 0, 20, 54, 61, 65, 72, 78, 85, 94, 104, 114, 121, 128, 132, 135, 136, 135, 132, 127, 120, 113, 110, 74, 6, 0, 0, 0, 0 ),
		( 0, 0, 0, 0, 22, 62, 67, 71, 78, 85, 92, 99, 106, 116, 127, 135, 142, 148, 151, 152, 151, 148, 141, 134, 125, 114, 109, 73, 3, 0, 0, 0 ),
		( 0, 0, 0, 18, 68, 73, 77, 83, 90, 97, 105, 112, 121, 128, 138, 148, 156, 163, 167, 168, 167, 162, 155, 147, 137, 126, 114, 108, 58, 0, 0, 0 ),
		( 0, 0, 7, 70, 80, 82, 88, 94, 101, 108, 116, 125, 133, 142, 151, 160, 171, 177, 182, 183, 181, 176, 169, 159, 148, 136, 123, 110, 100, 29, 0, 0 ),
		( 0, 0, 56, 90, 86, 91, 97, 103, 110, 118, 126, 135, 144, 153, 163, 172, 183, 191, 197, 199, 196, 190, 181, 170, 158, 145, 131, 116, 105, 80, 3, 0 ),
		( 0, 19, 99, 92, 95, 99, 105, 111, 118, 126, 134, 143, 153, 163, 174, 184, 195, 205, 213, 215, 211, 203, 192, 179, 166, 152, 137, 122, 107, 98, 31, 0 ),
		( 0, 65, 110, 99, 103, 106, 111, 118, 124, 132, 141, 150, 160, 170, 181, 193, 205, 217, 227, 231, 226, 214, 201, 186, 172, 157, 142, 126, 111, 99, 62, 0 ),
		( 13, 104, 113, 106, 109, 113, 118, 124, 130, 138, 145, 155, 165, 175, 186, 198, 212, 225, 239, 248, 237, 222, 206, 190, 175, 160, 143, 127, 112, 97, 78, 17 ),
		( 52, 125, 116, 112, 115, 119, 124, 129, 135, 142, 149, 158, 168, 178, 189, 200, 213, 226, 241, 249, 238, 222, 206, 190, 175, 160, 144, 128, 113, 96, 81, 38 ),
		( 94, 131, 122, 118, 122, 124, 129, 134, 139, 144, 152, 160, 169, 178, 188, 199, 210, 221, 230, 234, 228, 215, 202, 187, 172, 157, 142, 126, 111, 95, 78, 54 ),
		( 133, 136, 128, 124, 126, 129, 132, 136, 141, 147, 153, 161, 169, 176, 185, 194, 204, 212, 218, 219, 215, 205, 193, 180, 167, 152, 138, 122, 107, 92, 75, 63 ),
		( 151, 144, 136, 130, 131, 133, 135, 140, 143, 148, 154, 161, 167, 174, 181, 189, 196, 202, 206, 206, 202, 194, 183, 171, 159, 145, 131, 117, 103, 88, 71, 59 ),
		( 156, 150, 143, 136, 135, 136, 139, 142, 145, 149, 154, 159, 165, 171, 176, 183, 188, 191, 194, 193, 190, 183, 174, 162, 149, 137, 124, 111, 97, 82, 66, 54 ),
		( 165, 157, 150, 143, 139, 140, 141, 144, 147, 150, 153, 157, 162, 167, 171, 175, 179, 182, 183, 182, 179, 172, 163, 153, 139, 127, 115, 102, 88, 75, 60, 48 ),
		( 160, 164, 156, 150, 144, 143, 144, 145, 148, 150, 153, 155, 159, 163, 166, 169, 171, 173, 173, 171, 167, 162, 153, 143, 131, 118, 105, 93, 80, 68, 53, 34 ),
		( 125, 172, 163, 156, 150, 147, 147, 147, 148, 150, 151, 154, 156, 158, 161, 163, 164, 165, 163, 161, 157, 152, 144, 134, 123, 110, 96, 82, 71, 59, 45, 19 ),
		( 78, 181, 170, 164, 157, 151, 149, 149, 149, 149, 151, 152, 153, 155, 156, 157, 157, 157, 155, 152, 148, 142, 134, 126, 115, 103, 90, 74, 61, 49, 35, 6 ),
		( 23, 167, 182, 170, 164, 157, 152, 152, 150, 150, 150, 151, 151, 151, 151, 152, 150, 149, 147, 144, 140, 133, 126, 118, 107, 96, 83, 68, 53, 39, 21, 0 ),
		( 0, 119, 197, 176, 170, 163, 157, 153, 152, 151, 150, 149, 149, 149, 148, 146, 146, 143, 140, 136, 131, 126, 118, 109, 100, 88, 76, 62, 47, 31, 7, 0 ),
		( 0, 42, 202, 185, 177, 170, 163, 156, 153, 152, 150, 148, 147, 146, 145, 143, 140, 138, 134, 130, 124, 119, 111, 102, 93, 82, 70, 56, 42, 25, 0, 0 ),
		( 0, 0, 133, 206, 183, 177, 170, 163, 157, 153, 150, 148, 146, 144, 142, 139, 137, 133, 129, 124, 118, 112, 104, 96, 86, 76, 64, 51, 37, 13, 0, 0 ),
		( 0, 0, 25, 188, 198, 184, 177, 171, 164, 157, 151, 149, 146, 143, 140, 136, 133, 129, 124, 119, 113, 107, 99, 90, 81, 71, 58, 47, 30, 2, 0, 0 ),
		( 0, 0, 0, 64, 208, 195, 184, 177, 170, 164, 157, 151, 146, 142, 139, 135, 130, 126, 121, 115, 108, 102, 94, 85, 75, 64, 54, 46, 11, 0, 0, 0 ),
		( 0, 0, 0, 0, 87, 210, 196, 184, 177, 171, 164, 157, 150, 144, 139, 133, 129, 124, 118, 112, 105, 98, 90, 80, 71, 65, 60, 21, 0, 0, 0, 0 ),
		( 0, 0, 0, 0, 0, 81, 201, 202, 183, 177, 171, 164, 157, 151, 144, 137, 130, 124, 117, 111, 104, 97, 91, 84, 82, 72, 25, 0, 0, 0, 0, 0 ),
		( 0, 0, 0, 0, 0, 0, 49, 168, 207, 192, 177, 170, 164, 157, 151, 144, 137, 130, 124, 117, 111, 104, 101, 99, 71, 18, 0, 0, 0, 0, 0, 0 ),
		( 0, 0, 0, 0, 0, 0, 0, 6, 94, 164, 189, 179, 172, 165, 158, 151, 145, 138, 131, 125, 119, 113, 89, 46, 2, 0, 0, 0, 0, 0, 0, 0 ),
		( 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 94, 174, 181, 171, 164, 157, 151, 144, 137, 133, 117, 58, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0 )
	);
	
	
	constant WALL_SIZE_40 : integer := 40;
	type WALL40_COLOR_TYPE is array ( 0 to WALL_SIZE_40 - 1, 0 to  WALL_SIZE_40 - 1 ) of integer;
	constant WALL40_COLOR_R : WALL40_COLOR_TYPE := (
		( 107, 109, 112, 93, 85, 104, 117, 90, 91, 92, 89, 92, 115, 89, 77, 84, 88, 90, 83, 98, 98, 100, 114, 100, 87, 93, 110, 89, 84, 96, 90, 81, 88, 89, 93, 91, 94, 102, 94, 105 ),
		( 107, 111, 115, 95, 87, 104, 116, 92, 85, 87, 90, 90, 115, 86, 79, 85, 81, 91, 84, 101, 100, 100, 114, 100, 86, 93, 117, 90, 81, 95, 86, 80, 89, 87, 93, 83, 96, 100, 92, 104 ),
		( 110, 111, 116, 95, 83, 101, 118, 98, 90, 84, 91, 88, 115, 84, 78, 89, 79, 94, 89, 102, 98, 101, 114, 97, 88, 94, 118, 95, 83, 97, 87, 78, 84, 85, 92, 88, 95, 97, 94, 100 ),
		( 109, 111, 116, 97, 86, 104, 119, 103, 87, 82, 90, 85, 117, 91, 77, 87, 84, 91, 89, 100, 99, 102, 114, 98, 90, 93, 116, 95, 90, 94, 82, 75, 81, 84, 88, 85, 91, 94, 94, 97 ),
		( 108, 111, 117, 101, 89, 104, 120, 104, 88, 86, 90, 88, 116, 89, 80, 87, 84, 82, 78, 102, 102, 105, 113, 99, 91, 93, 115, 98, 79, 89, 85, 76, 91, 92, 87, 86, 90, 93, 94, 96 ),
		( 107, 110, 114, 103, 94, 105, 114, 104, 87, 86, 86, 85, 115, 81, 77, 88, 87, 83, 73, 104, 104, 106, 113, 102, 91, 90, 111, 96, 76, 83, 87, 79, 92, 91, 91, 87, 89, 90, 93, 94 ),
		( 107, 112, 111, 106, 93, 105, 113, 102, 80, 91, 82, 81, 115, 82, 75, 92, 93, 86, 78, 106, 106, 106, 113, 101, 92, 94, 110, 93, 79, 84, 92, 82, 94, 95, 93, 84, 87, 89, 89, 94 ),
		( 109, 112, 109, 108, 95, 107, 112, 99, 82, 89, 79, 82, 112, 80, 71, 94, 89, 86, 83, 107, 107, 108, 113, 102, 94, 91, 108, 90, 77, 91, 96, 78, 94, 93, 92, 84, 81, 84, 87, 98 ),
		( 110, 111, 106, 109, 99, 108, 109, 98, 83, 87, 79, 82, 106, 83, 81, 93, 91, 85, 90, 111, 113, 108, 111, 103, 92, 87, 105, 83, 77, 91, 93, 79, 90, 90, 88, 80, 84, 77, 74, 102 ),
		( 110, 112, 106, 107, 100, 107, 105, 96, 87, 93, 83, 82, 103, 79, 83, 95, 94, 87, 86, 110, 114, 110, 110, 102, 96, 85, 100, 81, 74, 89, 90, 77, 95, 94, 88, 83, 85, 79, 74, 99 ),
		( 108, 112, 104, 101, 105, 108, 103, 96, 87, 93, 86, 83, 100, 87, 83, 89, 87, 79, 85, 111, 113, 115, 112, 99, 94, 88, 97, 84, 78, 80, 87, 82, 98, 90, 82, 79, 80, 79, 81, 95 ),
		( 108, 112, 102, 99, 106, 106, 100, 85, 89, 89, 92, 86, 102, 88, 82, 91, 88, 84, 81, 107, 116, 117, 111, 99, 95, 92, 97, 84, 75, 77, 92, 81, 92, 88, 86, 82, 81, 79, 79, 98 ),
		( 107, 112, 101, 98, 106, 108, 98, 83, 87, 87, 90, 91, 100, 96, 89, 88, 93, 85, 77, 103, 116, 115, 111, 103, 97, 87, 99, 85, 80, 83, 90, 82, 92, 93, 89, 81, 80, 81, 83, 101 ),
		( 107, 110, 104, 97, 104, 110, 92, 81, 89, 90, 93, 91, 100, 91, 88, 87, 91, 88, 76, 100, 116, 114, 111, 101, 94, 89, 102, 91, 83, 83, 93, 86, 95, 92, 88, 84, 79, 88, 86, 101 ),
		( 108, 113, 105, 98, 104, 110, 89, 77, 89, 88, 94, 88, 99, 95, 88, 84, 90, 88, 77, 99, 113, 114, 111, 99, 90, 91, 102, 87, 86, 86, 94, 88, 92, 91, 92, 85, 72, 92, 92, 101 ),
		( 109, 114, 106, 95, 104, 114, 90, 80, 87, 90, 87, 97, 102, 93, 82, 87, 94, 88, 76, 96, 110, 115, 107, 97, 89, 95, 104, 84, 89, 90, 90, 90, 88, 93, 94, 84, 76, 93, 88, 101 ),
		( 107, 114, 104, 92, 104, 115, 92, 77, 90, 92, 88, 90, 102, 86, 84, 89, 95, 88, 79, 96, 109, 113, 108, 95, 89, 92, 108, 81, 85, 83, 79, 88, 90, 96, 95, 86, 74, 94, 94, 103 ),
		( 108, 113, 104, 94, 102, 116, 91, 78, 91, 90, 83, 95, 101, 83, 81, 92, 95, 89, 79, 93, 106, 113, 110, 95, 86, 92, 105, 86, 89, 84, 83, 86, 82, 96, 98, 93, 72, 91, 90, 104 ),
		( 106, 113, 102, 85, 97, 118, 94, 76, 87, 89, 81, 100, 100, 77, 80, 89, 89, 82, 81, 95, 106, 114, 108, 97, 87, 93, 106, 87, 88, 77, 87, 85, 80, 91, 96, 92, 77, 88, 89, 107 ),
		( 105, 112, 99, 83, 95, 119, 96, 76, 83, 87, 86, 97, 100, 76, 76, 89, 94, 85, 76, 94, 105, 114, 109, 97, 88, 93, 105, 86, 90, 80, 89, 85, 80, 94, 96, 87, 76, 84, 79, 111 ),
		( 102, 111, 94, 84, 98, 119, 98, 79, 87, 89, 83, 95, 101, 76, 79, 83, 91, 89, 73, 94, 101, 115, 110, 95, 86, 95, 97, 88, 98, 85, 86, 86, 88, 96, 95, 88, 83, 80, 84, 113 ),
		( 100, 109, 98, 83, 97, 118, 95, 72, 89, 92, 82, 97, 100, 73, 80, 86, 93, 88, 72, 90, 100, 113, 109, 93, 86, 99, 94, 88, 94, 91, 87, 88, 85, 92, 92, 86, 84, 80, 83, 113 ),
		( 97, 113, 97, 82, 95, 117, 94, 72, 80, 89, 88, 97, 104, 73, 82, 84, 95, 89, 74, 91, 101, 112, 109, 92, 86, 101, 94, 88, 91, 90, 86, 88, 85, 92, 92, 90, 90, 82, 86, 114 ),
		( 96, 113, 99, 86, 95, 117, 97, 80, 81, 87, 93, 93, 102, 73, 91, 90, 91, 87, 74, 85, 99, 113, 110, 95, 86, 95, 94, 82, 88, 93, 88, 91, 86, 89, 94, 93, 85, 81, 87, 113 ),
		( 96, 112, 101, 86, 93, 118, 96, 78, 86, 86, 91, 93, 105, 82, 91, 89, 86, 86, 79, 85, 95, 111, 105, 93, 87, 98, 95, 81, 83, 91, 89, 95, 89, 88, 92, 93, 92, 82, 93, 114 ),
		( 95, 112, 101, 88, 93, 116, 94, 76, 89, 87, 94, 96, 103, 84, 86, 89, 86, 86, 80, 83, 95, 114, 106, 92, 85, 97, 96, 83, 87, 93, 93, 90, 89, 89, 89, 95, 93, 82, 97, 115 ),
		( 99, 111, 105, 88, 91, 114, 95, 80, 93, 88, 94, 96, 102, 81, 89, 92, 87, 87, 72, 80, 91, 115, 106, 95, 88, 94, 99, 84, 80, 88, 94, 87, 83, 87, 88, 85, 96, 85, 100, 113 ),
		( 98, 109, 105, 89, 90, 114, 98, 85, 93, 83, 91, 99, 104, 82, 86, 87, 83, 86, 79, 79, 91, 116, 106, 95, 91, 100, 97, 83, 79, 84, 96, 90, 87, 88, 86, 85, 96, 89, 106, 110 ),
		( 96, 109, 105, 86, 87, 112, 96, 84, 88, 81, 90, 103, 106, 83, 81, 84, 83, 86, 77, 80, 94, 113, 106, 97, 87, 99, 97, 77, 82, 83, 97, 89, 87, 85, 84, 90, 96, 90, 108, 108 ),
		( 96, 106, 105, 89, 86, 110, 99, 86, 91, 82, 88, 105, 107, 86, 85, 84, 87, 82, 78, 83, 95, 106, 104, 98, 88, 101, 93, 79, 85, 87, 103, 89, 90, 83, 87, 97, 93, 96, 110, 103 ),
		( 97, 106, 107, 89, 87, 105, 103, 83, 89, 77, 87, 105, 109, 90, 88, 82, 89, 86, 73, 86, 94, 105, 105, 95, 86, 98, 93, 77, 89, 94, 104, 95, 98, 84, 88, 95, 86, 99, 112, 100 ),
		( 99, 107, 105, 95, 90, 106, 102, 81, 86, 80, 83, 110, 113, 91, 84, 78, 93, 88, 74, 85, 95, 105, 106, 93, 93, 97, 96, 76, 90, 101, 104, 92, 89, 84, 92, 83, 89, 104, 111, 105 ),
		( 99, 107, 105, 91, 88, 102, 107, 80, 86, 85, 76, 113, 115, 94, 82, 79, 90, 88, 82, 82, 91, 105, 110, 93, 90, 99, 100, 80, 94, 102, 106, 88, 92, 87, 92, 81, 87, 113, 110, 109 ),
		( 101, 108, 108, 90, 88, 102, 111, 85, 80, 83, 80, 108, 118, 94, 81, 84, 96, 84, 81, 84, 92, 104, 110, 94, 88, 99, 101, 89, 88, 96, 110, 89, 86, 84, 88, 85, 87, 114, 109, 107 ),
		( 101, 106, 110, 89, 86, 103, 113, 91, 86, 88, 81, 109, 118, 92, 78, 85, 90, 83, 91, 86, 92, 106, 110, 95, 90, 93, 102, 88, 79, 95, 114, 88, 89, 89, 85, 86, 92, 114, 111, 109 ),
		( 104, 107, 113, 93, 86, 104, 115, 89, 84, 95, 81, 107, 116, 96, 82, 83, 83, 85, 92, 88, 95, 107, 112, 97, 96, 94, 99, 87, 79, 94, 114, 89, 88, 87, 85, 88, 92, 116, 113, 110 ),
		( 104, 108, 112, 95, 87, 106, 117, 87, 78, 96, 83, 105, 117, 89, 80, 85, 85, 87, 94, 91, 93, 106, 112, 97, 94, 95, 99, 89, 80, 95, 112, 86, 86, 93, 85, 87, 89, 116, 110, 108 ),
		( 105, 108, 113, 95, 92, 105, 117, 94, 84, 92, 92, 100, 114, 94, 84, 88, 80, 89, 93, 92, 97, 104, 115, 100, 97, 95, 100, 92, 82, 93, 105, 83, 86, 93, 93, 82, 90, 113, 102, 109 ),
		( 105, 109, 112, 96, 90, 102, 116, 91, 88, 90, 89, 96, 114, 92, 81, 87, 76, 82, 85, 91, 101, 103, 113, 99, 96, 95, 102, 92, 77, 92, 98, 86, 89, 90, 92, 85, 93, 109, 97, 111 ),
		( 107, 111, 113, 96, 90, 103, 117, 93, 86, 87, 86, 95, 115, 94, 78, 87, 81, 87, 84, 95, 100, 102, 113, 100, 93, 97, 107, 91, 76, 91, 94, 89, 89, 89, 96, 87, 96, 103, 95, 112 )
	);
	constant WALL40_COLOR_G : WALL40_COLOR_TYPE := (
		( 66, 68, 69, 54, 49, 63, 72, 52, 53, 55, 52, 54, 70, 53, 45, 50, 52, 54, 49, 58, 59, 59, 70, 59, 50, 56, 67, 51, 47, 56, 51, 46, 53, 53, 55, 55, 55, 61, 55, 64 ),
		( 66, 68, 71, 56, 51, 62, 72, 53, 49, 51, 52, 53, 70, 50, 46, 51, 47, 55, 49, 60, 59, 59, 70, 59, 49, 55, 72, 52, 46, 56, 48, 46, 54, 50, 55, 49, 56, 60, 53, 61 ),
		( 67, 68, 71, 56, 48, 61, 72, 58, 52, 49, 52, 51, 71, 49, 46, 52, 46, 56, 52, 60, 58, 60, 70, 57, 51, 56, 73, 56, 47, 57, 49, 44, 50, 49, 55, 52, 55, 57, 55, 59 ),
		( 67, 68, 70, 58, 51, 62, 73, 62, 50, 48, 53, 49, 71, 52, 44, 52, 50, 54, 52, 60, 59, 61, 70, 58, 52, 55, 72, 56, 52, 55, 46, 43, 48, 49, 53, 52, 53, 55, 55, 58 ),
		( 67, 68, 72, 61, 52, 63, 74, 63, 51, 50, 52, 50, 71, 52, 46, 52, 50, 49, 44, 60, 62, 63, 69, 59, 53, 55, 71, 57, 46, 51, 48, 44, 54, 54, 52, 50, 53, 54, 55, 57 ),
		( 65, 68, 69, 62, 56, 63, 70, 62, 50, 51, 49, 49, 71, 47, 44, 52, 50, 49, 42, 62, 63, 64, 69, 61, 53, 53, 68, 57, 44, 47, 50, 45, 55, 53, 54, 51, 52, 52, 54, 56 ),
		( 65, 69, 67, 64, 55, 63, 69, 60, 45, 54, 47, 46, 70, 47, 43, 56, 55, 51, 45, 64, 63, 64, 69, 61, 53, 56, 67, 55, 46, 47, 53, 47, 56, 56, 55, 50, 51, 51, 52, 55 ),
		( 66, 68, 66, 66, 56, 64, 68, 59, 47, 52, 44, 47, 68, 45, 41, 58, 53, 51, 48, 64, 64, 65, 70, 61, 54, 53, 65, 53, 44, 52, 56, 45, 56, 55, 55, 50, 47, 49, 50, 57 ),
		( 66, 68, 64, 66, 59, 65, 66, 58, 48, 51, 45, 47, 64, 47, 48, 58, 54, 50, 53, 67, 69, 65, 68, 61, 54, 50, 63, 49, 45, 53, 55, 46, 53, 53, 52, 48, 48, 44, 42, 59 ),
		( 67, 69, 64, 65, 59, 64, 63, 57, 50, 55, 48, 46, 62, 45, 49, 58, 56, 51, 49, 67, 70, 66, 68, 61, 57, 49, 59, 47, 43, 53, 53, 44, 56, 55, 52, 50, 49, 45, 42, 57 ),
		( 65, 68, 62, 61, 62, 65, 61, 57, 51, 55, 51, 47, 60, 50, 49, 53, 52, 47, 49, 68, 69, 70, 69, 59, 55, 51, 57, 49, 46, 48, 51, 46, 59, 53, 48, 47, 46, 46, 47, 56 ),
		( 66, 69, 61, 59, 64, 64, 59, 49, 51, 52, 54, 50, 61, 51, 48, 55, 53, 50, 46, 65, 72, 72, 68, 60, 55, 53, 57, 49, 44, 44, 55, 46, 55, 53, 51, 48, 46, 46, 46, 58 ),
		( 65, 69, 60, 58, 64, 65, 58, 48, 51, 50, 53, 52, 59, 55, 53, 53, 55, 50, 43, 63, 71, 71, 69, 62, 56, 51, 59, 50, 47, 49, 55, 46, 55, 55, 52, 48, 45, 47, 48, 59 ),
		( 66, 67, 63, 58, 63, 67, 54, 46, 52, 52, 54, 52, 59, 53, 53, 52, 55, 52, 42, 59, 71, 70, 68, 61, 54, 52, 61, 53, 48, 49, 56, 49, 57, 55, 51, 49, 45, 52, 50, 60 ),
		( 66, 69, 63, 58, 63, 67, 52, 44, 51, 50, 54, 50, 59, 56, 53, 49, 54, 51, 43, 59, 69, 70, 68, 59, 52, 53, 60, 51, 51, 51, 57, 50, 55, 54, 53, 50, 41, 54, 54, 61 ),
		( 66, 70, 64, 55, 63, 70, 53, 46, 50, 52, 50, 56, 60, 54, 48, 51, 57, 52, 42, 58, 66, 70, 65, 57, 51, 56, 62, 50, 53, 54, 53, 52, 52, 55, 55, 50, 44, 55, 51, 60 ),
		( 65, 70, 62, 54, 63, 71, 53, 43, 52, 53, 51, 52, 60, 50, 50, 52, 57, 51, 45, 57, 66, 69, 67, 57, 51, 54, 65, 48, 51, 49, 46, 51, 54, 58, 56, 51, 43, 55, 55, 61 ),
		( 66, 69, 62, 54, 62, 72, 53, 44, 52, 51, 48, 55, 60, 48, 48, 54, 56, 52, 45, 54, 64, 70, 68, 56, 50, 53, 62, 51, 53, 50, 49, 49, 47, 57, 58, 56, 41, 54, 53, 63 ),
		( 64, 69, 61, 50, 58, 72, 54, 43, 50, 51, 46, 58, 58, 44, 47, 52, 52, 48, 47, 55, 64, 69, 67, 57, 50, 54, 63, 51, 53, 46, 52, 47, 46, 55, 57, 55, 44, 52, 52, 64 ),
		( 64, 68, 59, 48, 57, 72, 56, 43, 47, 50, 49, 57, 59, 43, 45, 53, 55, 51, 43, 55, 63, 70, 67, 58, 51, 55, 62, 52, 55, 47, 53, 48, 46, 57, 57, 51, 43, 49, 46, 67 ),
		( 62, 68, 55, 48, 58, 72, 58, 46, 49, 52, 47, 56, 60, 43, 47, 49, 53, 53, 41, 56, 60, 70, 68, 56, 49, 56, 57, 52, 59, 51, 51, 48, 51, 57, 56, 52, 47, 45, 49, 69 ),
		( 60, 67, 57, 48, 57, 71, 56, 40, 51, 54, 47, 58, 60, 42, 47, 49, 54, 52, 40, 52, 60, 69, 67, 55, 49, 59, 56, 51, 56, 55, 51, 50, 49, 55, 55, 51, 47, 46, 47, 69 ),
		( 58, 69, 58, 47, 56, 71, 55, 40, 46, 52, 51, 57, 62, 41, 48, 49, 56, 54, 42, 53, 60, 69, 66, 54, 50, 60, 55, 52, 53, 53, 50, 49, 49, 55, 54, 52, 52, 46, 50, 69 ),
		( 57, 69, 60, 50, 56, 71, 56, 46, 47, 50, 54, 55, 61, 41, 54, 53, 54, 53, 43, 49, 58, 69, 67, 55, 49, 56, 55, 47, 51, 55, 51, 53, 50, 53, 56, 55, 49, 45, 51, 69 ),
		( 57, 69, 60, 50, 54, 72, 56, 44, 50, 49, 53, 54, 62, 48, 53, 52, 50, 51, 46, 48, 56, 67, 64, 55, 50, 58, 55, 47, 48, 54, 52, 55, 52, 53, 55, 56, 54, 46, 55, 70 ),
		( 56, 69, 60, 51, 55, 72, 55, 43, 52, 51, 56, 57, 61, 49, 50, 52, 50, 51, 46, 48, 56, 70, 65, 54, 49, 58, 57, 49, 50, 54, 54, 53, 53, 54, 53, 57, 54, 46, 58, 70 ),
		( 58, 68, 62, 51, 53, 70, 57, 46, 55, 51, 55, 57, 61, 47, 53, 54, 50, 52, 41, 45, 53, 71, 65, 55, 51, 56, 58, 48, 46, 51, 55, 50, 50, 52, 52, 50, 56, 49, 60, 69 ),
		( 57, 66, 63, 51, 53, 69, 58, 49, 55, 48, 53, 59, 62, 47, 51, 50, 48, 51, 45, 45, 53, 71, 64, 55, 53, 60, 57, 48, 46, 49, 56, 51, 52, 53, 51, 50, 56, 51, 64, 67 ),
		( 56, 66, 64, 50, 51, 69, 56, 49, 52, 46, 52, 61, 64, 47, 48, 49, 48, 50, 44, 45, 55, 69, 64, 57, 51, 59, 57, 44, 47, 48, 57, 50, 52, 51, 49, 54, 57, 53, 66, 64 ),
		( 57, 65, 63, 52, 49, 67, 59, 49, 54, 47, 51, 63, 64, 49, 51, 49, 51, 48, 44, 48, 56, 64, 63, 57, 51, 60, 54, 45, 49, 51, 62, 51, 54, 49, 51, 58, 54, 56, 67, 62 ),
		( 57, 64, 64, 51, 50, 63, 62, 48, 53, 44, 50, 63, 66, 52, 53, 48, 51, 51, 42, 50, 55, 63, 64, 55, 49, 58, 54, 43, 51, 55, 62, 55, 59, 49, 52, 57, 50, 59, 68, 59 ),
		( 58, 65, 63, 55, 52, 64, 61, 46, 50, 46, 47, 66, 68, 53, 50, 45, 54, 52, 44, 49, 55, 63, 64, 54, 54, 58, 57, 43, 52, 60, 62, 54, 53, 49, 55, 49, 52, 63, 67, 63 ),
		( 59, 65, 64, 53, 51, 62, 65, 46, 51, 49, 42, 69, 71, 55, 48, 46, 52, 52, 48, 47, 53, 64, 66, 54, 52, 60, 59, 45, 55, 61, 64, 51, 56, 51, 55, 46, 51, 69, 68, 67 ),
		( 61, 66, 66, 52, 51, 62, 66, 49, 48, 48, 45, 66, 73, 55, 48, 49, 56, 50, 48, 49, 54, 62, 67, 55, 51, 59, 60, 51, 52, 57, 67, 52, 52, 50, 53, 49, 50, 69, 66, 66 ),
		( 61, 65, 66, 52, 49, 61, 68, 54, 51, 53, 46, 67, 72, 54, 46, 50, 52, 49, 53, 50, 54, 64, 68, 55, 52, 55, 60, 50, 45, 56, 70, 51, 53, 53, 51, 49, 53, 70, 68, 66 ),
		( 62, 65, 69, 55, 49, 62, 71, 52, 51, 57, 47, 65, 71, 56, 49, 49, 48, 50, 55, 51, 56, 65, 69, 56, 56, 56, 59, 51, 45, 55, 70, 51, 53, 51, 50, 51, 53, 70, 68, 66 ),
		( 62, 66, 68, 56, 50, 64, 71, 50, 47, 58, 48, 64, 72, 52, 47, 50, 49, 51, 56, 52, 55, 64, 69, 57, 55, 57, 60, 51, 45, 56, 68, 49, 52, 55, 51, 50, 52, 71, 67, 65 ),
		( 64, 66, 69, 56, 53, 64, 72, 54, 49, 56, 53, 60, 70, 55, 50, 52, 46, 53, 54, 54, 57, 62, 70, 59, 56, 56, 59, 54, 47, 54, 63, 48, 51, 55, 56, 47, 53, 68, 61, 66 ),
		( 64, 67, 69, 57, 52, 61, 71, 53, 52, 55, 52, 57, 70, 54, 48, 51, 43, 49, 50, 53, 60, 62, 70, 58, 56, 56, 61, 54, 43, 54, 58, 50, 53, 53, 56, 50, 54, 66, 57, 68 ),
		( 66, 69, 70, 57, 52, 61, 72, 53, 50, 52, 49, 55, 70, 56, 46, 52, 46, 52, 49, 55, 59, 62, 70, 60, 54, 58, 65, 52, 43, 53, 55, 51, 54, 52, 57, 52, 56, 62, 56, 69 )
	);
	constant WALL40_COLOR_B : WALL40_COLOR_TYPE := (
		( 37, 39, 39, 32, 29, 35, 41, 31, 32, 33, 30, 32, 40, 30, 28, 31, 31, 32, 29, 33, 34, 34, 39, 33, 29, 33, 38, 31, 27, 32, 30, 28, 32, 31, 34, 32, 31, 34, 32, 36 ),
		( 38, 39, 39, 32, 30, 35, 40, 31, 29, 33, 30, 30, 39, 28, 28, 31, 29, 33, 29, 34, 35, 35, 40, 33, 29, 32, 41, 30, 26, 32, 29, 27, 33, 30, 33, 30, 31, 33, 31, 35 ),
		( 40, 39, 40, 32, 29, 34, 41, 33, 30, 31, 31, 30, 40, 28, 28, 32, 28, 34, 30, 34, 33, 34, 39, 33, 30, 33, 41, 32, 27, 32, 29, 27, 31, 29, 32, 31, 31, 32, 32, 34 ),
		( 39, 39, 39, 33, 30, 35, 41, 35, 29, 30, 30, 29, 41, 30, 27, 32, 30, 33, 30, 34, 34, 34, 40, 34, 30, 32, 40, 32, 30, 31, 27, 26, 29, 28, 32, 30, 31, 31, 31, 33 ),
		( 39, 39, 39, 34, 31, 35, 42, 36, 30, 32, 31, 30, 40, 30, 28, 32, 29, 30, 27, 35, 35, 36, 40, 33, 30, 31, 40, 33, 28, 29, 27, 26, 33, 32, 31, 30, 30, 30, 31, 33 ),
		( 38, 39, 38, 35, 32, 35, 39, 35, 29, 31, 30, 29, 40, 27, 28, 32, 30, 30, 26, 36, 35, 36, 40, 35, 31, 31, 39, 33, 27, 27, 29, 26, 33, 31, 32, 30, 30, 29, 31, 33 ),
		( 37, 39, 37, 37, 31, 35, 38, 34, 26, 32, 30, 27, 39, 28, 27, 34, 33, 32, 27, 36, 36, 36, 40, 34, 31, 32, 38, 31, 28, 27, 31, 27, 33, 33, 33, 30, 29, 29, 29, 32 ),
		( 37, 38, 37, 37, 33, 35, 38, 34, 27, 31, 28, 28, 37, 27, 26, 35, 32, 31, 28, 36, 37, 37, 40, 35, 31, 31, 37, 31, 27, 30, 32, 27, 34, 33, 33, 30, 27, 27, 28, 33 ),
		( 37, 38, 36, 36, 34, 36, 37, 34, 28, 30, 28, 28, 36, 28, 30, 35, 34, 31, 30, 37, 38, 37, 39, 35, 30, 29, 36, 29, 28, 30, 33, 27, 32, 32, 31, 29, 28, 24, 24, 34 ),
		( 37, 39, 36, 37, 34, 37, 36, 33, 29, 31, 29, 27, 35, 27, 30, 35, 34, 31, 29, 36, 39, 37, 39, 34, 32, 28, 33, 28, 27, 31, 32, 26, 34, 33, 31, 30, 28, 25, 24, 32 ),
		( 37, 39, 35, 35, 35, 37, 35, 32, 29, 31, 30, 28, 34, 30, 30, 32, 32, 29, 28, 37, 39, 39, 40, 34, 31, 29, 33, 29, 27, 29, 32, 27, 35, 31, 29, 29, 27, 26, 27, 32 ),
		( 37, 39, 34, 34, 36, 36, 34, 29, 30, 28, 31, 28, 34, 30, 30, 33, 32, 30, 27, 36, 40, 40, 40, 34, 31, 31, 32, 28, 26, 27, 33, 27, 33, 31, 30, 30, 28, 28, 27, 33 ),
		( 37, 39, 35, 34, 36, 36, 33, 27, 30, 28, 30, 30, 34, 33, 32, 32, 33, 30, 26, 36, 40, 40, 39, 35, 31, 29, 33, 29, 27, 29, 32, 27, 32, 33, 31, 30, 27, 28, 28, 34 ),
		( 37, 37, 35, 33, 36, 38, 32, 28, 31, 29, 31, 30, 34, 31, 32, 32, 33, 30, 26, 33, 39, 39, 39, 34, 31, 30, 34, 31, 28, 30, 34, 28, 33, 32, 31, 30, 27, 30, 28, 34 ),
		( 38, 39, 36, 33, 36, 37, 31, 26, 30, 29, 29, 29, 33, 32, 32, 30, 33, 30, 25, 33, 38, 39, 40, 34, 30, 31, 34, 30, 30, 31, 33, 29, 32, 33, 31, 30, 25, 32, 30, 35 ),
		( 37, 39, 36, 32, 35, 38, 31, 26, 29, 30, 28, 32, 35, 32, 30, 31, 34, 31, 25, 34, 37, 39, 37, 33, 30, 32, 34, 30, 33, 33, 32, 30, 30, 33, 32, 31, 25, 31, 28, 34 ),
		( 38, 40, 36, 31, 36, 39, 31, 26, 30, 31, 29, 30, 34, 29, 31, 31, 34, 31, 27, 33, 37, 38, 38, 32, 29, 31, 35, 28, 32, 31, 28, 28, 31, 34, 33, 31, 25, 32, 30, 35 ),
		( 39, 40, 35, 32, 35, 40, 31, 26, 30, 30, 27, 31, 33, 28, 29, 31, 32, 32, 26, 32, 36, 39, 40, 32, 28, 31, 34, 30, 33, 32, 29, 28, 30, 34, 34, 33, 25, 31, 29, 35 ),
		( 37, 39, 35, 29, 34, 40, 32, 25, 28, 30, 26, 33, 33, 26, 29, 30, 31, 30, 27, 32, 36, 39, 39, 33, 29, 31, 34, 32, 32, 29, 30, 28, 29, 33, 34, 33, 26, 29, 29, 36 ),
		( 37, 39, 33, 29, 33, 40, 32, 25, 27, 29, 28, 32, 33, 26, 28, 30, 32, 31, 26, 33, 35, 39, 39, 33, 29, 32, 35, 31, 32, 29, 30, 28, 28, 34, 34, 31, 26, 28, 27, 38 ),
		( 35, 38, 32, 28, 33, 39, 33, 27, 28, 30, 28, 31, 34, 26, 30, 29, 31, 33, 25, 32, 34, 39, 40, 33, 29, 32, 32, 31, 34, 31, 29, 28, 30, 34, 33, 32, 27, 26, 28, 39 ),
		( 35, 38, 33, 28, 33, 39, 32, 24, 29, 31, 28, 33, 34, 26, 30, 29, 32, 33, 25, 30, 33, 39, 39, 32, 28, 33, 32, 30, 32, 33, 30, 29, 29, 33, 32, 32, 28, 26, 28, 40 ),
		( 34, 39, 33, 28, 32, 39, 31, 24, 26, 30, 30, 32, 35, 26, 31, 29, 33, 33, 25, 30, 34, 39, 39, 30, 29, 34, 32, 31, 31, 32, 28, 30, 30, 33, 32, 32, 30, 26, 29, 39 ),
		( 33, 39, 34, 29, 32, 39, 32, 27, 27, 29, 31, 31, 35, 25, 32, 31, 31, 32, 26, 29, 33, 39, 39, 31, 29, 33, 31, 29, 30, 31, 29, 30, 30, 32, 34, 33, 28, 26, 29, 39 ),
		( 32, 39, 33, 29, 32, 40, 32, 26, 29, 28, 31, 31, 35, 28, 33, 30, 29, 32, 27, 28, 32, 38, 37, 31, 29, 33, 31, 28, 28, 30, 30, 32, 32, 32, 33, 33, 31, 27, 31, 40 ),
		( 31, 38, 34, 29, 32, 40, 32, 25, 31, 29, 32, 32, 35, 30, 32, 30, 29, 32, 28, 28, 32, 40, 37, 30, 28, 34, 32, 29, 29, 30, 31, 31, 32, 32, 32, 34, 31, 27, 32, 41 ),
		( 33, 39, 36, 30, 31, 39, 32, 27, 32, 29, 32, 32, 34, 28, 32, 31, 29, 32, 26, 27, 31, 39, 37, 31, 30, 33, 33, 28, 27, 28, 31, 29, 31, 32, 32, 30, 32, 28, 34, 40 ),
		( 33, 38, 36, 29, 30, 39, 33, 28, 32, 28, 31, 34, 35, 28, 32, 30, 29, 32, 29, 26, 31, 39, 37, 30, 30, 35, 33, 27, 26, 28, 32, 30, 31, 32, 32, 30, 32, 30, 36, 38 ),
		( 32, 38, 36, 29, 29, 39, 33, 28, 30, 27, 31, 35, 36, 29, 30, 30, 28, 31, 27, 27, 32, 39, 37, 31, 29, 35, 33, 25, 28, 28, 33, 30, 31, 31, 31, 32, 32, 30, 37, 36 ),
		( 32, 38, 36, 30, 29, 38, 34, 29, 32, 28, 29, 35, 36, 28, 31, 30, 29, 30, 27, 28, 32, 36, 36, 32, 29, 35, 31, 26, 29, 30, 35, 30, 33, 31, 32, 34, 31, 32, 38, 34 ),
		( 32, 37, 36, 30, 29, 36, 35, 28, 32, 26, 29, 36, 37, 30, 32, 29, 30, 31, 25, 28, 32, 35, 37, 30, 29, 34, 32, 25, 30, 32, 34, 32, 35, 30, 32, 32, 29, 33, 39, 34 ),
		( 33, 37, 36, 32, 30, 37, 35, 27, 31, 28, 28, 37, 38, 31, 31, 27, 31, 32, 26, 28, 32, 35, 37, 30, 31, 34, 33, 25, 30, 34, 36, 31, 32, 31, 35, 30, 30, 35, 38, 37 ),
		( 34, 38, 36, 30, 29, 35, 37, 27, 31, 30, 26, 39, 39, 31, 29, 27, 30, 32, 28, 27, 31, 36, 38, 30, 30, 35, 34, 27, 31, 34, 36, 30, 34, 31, 33, 28, 29, 38, 38, 39 ),
		( 34, 38, 37, 30, 30, 35, 37, 28, 29, 29, 27, 37, 40, 31, 29, 29, 31, 31, 28, 28, 31, 35, 39, 30, 30, 34, 35, 29, 29, 33, 37, 30, 32, 30, 31, 29, 28, 39, 37, 37 ),
		( 34, 37, 37, 30, 29, 35, 38, 30, 31, 32, 27, 38, 41, 31, 28, 30, 30, 31, 31, 29, 32, 36, 39, 32, 30, 32, 35, 29, 27, 32, 39, 30, 32, 31, 30, 29, 30, 39, 38, 37 ),
		( 35, 37, 39, 32, 29, 35, 39, 29, 30, 34, 27, 37, 40, 32, 30, 30, 28, 31, 31, 30, 32, 36, 39, 31, 32, 33, 34, 29, 27, 32, 39, 30, 32, 30, 30, 30, 30, 38, 37, 36 ),
		( 36, 39, 38, 32, 29, 36, 39, 28, 28, 34, 27, 37, 40, 30, 28, 30, 29, 31, 32, 30, 31, 36, 39, 31, 32, 33, 35, 31, 26, 32, 38, 29, 32, 33, 31, 30, 30, 38, 37, 36 ),
		( 38, 39, 39, 32, 31, 36, 40, 31, 29, 34, 30, 35, 41, 32, 29, 32, 27, 31, 31, 31, 33, 36, 40, 33, 33, 33, 34, 31, 27, 31, 36, 29, 31, 33, 34, 29, 30, 37, 33, 37 ),
		( 37, 39, 39, 34, 30, 35, 40, 31, 31, 33, 30, 33, 40, 31, 29, 32, 26, 31, 29, 31, 34, 36, 40, 32, 32, 33, 35, 32, 26, 30, 34, 29, 32, 31, 34, 30, 31, 36, 33, 38 ),
		( 38, 40, 39, 33, 31, 35, 41, 31, 30, 33, 29, 32, 39, 32, 29, 31, 28, 31, 29, 32, 34, 35, 40, 33, 32, 33, 37, 31, 25, 30, 32, 31, 33, 32, 34, 30, 32, 34, 32, 38 )
	);

--    signal rom_addr, rom_col: unsigned(0 to 2);
--    signal rom_bit: std_logic;
    -- x, y coordinates of the ball
--    signal ball_x_l : unsigned(OBJECT_SIZE-1 downto 0);
--    signal ball_y_t : unsigned(OBJECT_SIZE-1 downto 0);
--    signal ball_x_r : unsigned(OBJECT_SIZE-1 downto 0);
--    signal ball_y_b : unsigned(OBJECT_SIZE-1 downto 0);

    -- signals that holds the x, y coordinates
--    signal pix_x, pix_y: unsigned (OBJECT_SIZE-1 downto 0);

--    signal wall_on, box_on, square_ball_on, ball_on: std_logic;
--    signal wall_rgb, box_rgb, ball_rgb: std_logic_vector(23 downto 0);
	
	-- ---------------------------------------------------------------------
	-- ---------------------------------------------------------------------
	-- ADDED BY MAKKUS
    signal pixelX : unsigned( OBJECT_SIZE - 1 downto 0 );
    signal pixelY : unsigned( OBJECT_SIZE - 1 downto 0 );
	
--	signal varShake : unsigned( OBJECT_SIZE - 1 downto 0 );
	signal varAddress : unsigned( OBJECT_SIZE - 1 downto 0 );
	signal varValue : unsigned( OBJECT_SIZE - 1 downto 0 );
	
--	signal varAddressBack1 : unsigned( OBJECT_SIZE - 1 downto 0 );
--	signal varValueBack1 : unsigned( OBJECT_SIZE - 1 downto 0 );
	
--	signal varAddressBack2 : unsigned( OBJECT_SIZE - 1 downto 0 );
--	signal varValueBack2 : unsigned( OBJECT_SIZE - 1 downto 0 );
		
	constant BALL_COUNT : integer := 16;
	
    type BALL_ARR_UNSIGNED is array ( 0 to BALL_COUNT - 1 ) of unsigned( OBJECT_SIZE - 1 downto 0 );
    type BALL_ARR_VECTOR is array ( 0 to BALL_COUNT - 1 ) of std_logic_vector( 23 downto 0 );
    type BALL_ARR_LOGIC is array ( 0 to BALL_COUNT - 1 ) of std_logic;
	
	signal ballMinX : BALL_ARR_UNSIGNED;
	signal ballMinY : BALL_ARR_UNSIGNED;
	signal ballMaxX : BALL_ARR_UNSIGNED;
	signal ballMaxY : BALL_ARR_UNSIGNED;
	signal ballOn : BALL_ARR_LOGIC;
	
	constant addressMinX : BALL_ARR_UNSIGNED := (
		x"0000",
		x"0002",
		x"0004",
		x"0006",
		x"0008",
		x"000A",
		x"000C",
		x"000E",
		x"0010",
		x"0012",
		x"0014",
		x"0016",
		x"0018",
		x"001A",
		x"001C",
		x"001E"
	);
	
	constant addressMinY : BALL_ARR_UNSIGNED := (
		x"0001",
		x"0003",
		x"0005",
		x"0007",
		x"0009",
		x"000B",
		x"000D",
		x"000F",
		x"0011",
		x"0013",
		x"0015",
		x"0017",
		x"0019",
		x"001B",
		x"001D",
		x"001F"
	);
	
	constant ballRgb : BALL_ARR_VECTOR := (
		x"FFFFFF",
		x"771177",
		x"117777",
		x"0000FF",
		x"FFFF00",
		x"000000",
		x"771111",
		x"111177",
		x"FF00FF",
		x"BB7711",
		x"FF0000",
		x"888888",
		x"00FFFF",
		x"777711",
		x"00FF00",
		x"117711"
	);
	
	
	signal pixVecR : std_logic_vector( 15 downto 0 );
	signal pixVecG : std_logic_vector( 15 downto 0 );
	signal pixVecB : std_logic_vector( 15 downto 0 );
	
	signal pixelIsBackground : boolean := true;
	
	signal ballIdx : integer;
	signal cueballIdx : integer;
	
	signal romX : integer;
	signal romY : integer;
	signal ballR : integer;
	signal ballG : integer;
	signal ballB : integer;
	signal shadeR : integer;
	signal shadeG : integer;
	signal shadeB : integer;
	signal shadeA : integer;
	signal pixR : integer;
	signal pixG : integer;
	signal pixB : integer;
	
	------
	
	
	signal pixelIsBall : boolean := false;
	signal pixelIsWall : boolean := false;
	signal pixelIsHole : boolean := false;
	signal pixelIsTable : boolean := false;
	signal pixelIsCueball : boolean := false;
	
	
		
	constant HOLE_COUNT : integer := 16;
	
    type HOLE_ARR_UNSIGNED is array ( 0 to HOLE_COUNT - 1 ) of unsigned( OBJECT_SIZE - 1 downto 0 );
    type HOLE_ARR_VECTOR is array ( 0 to HOLE_COUNT - 1 ) of std_logic_vector( 23 downto 0 );
    type HOLE_ARR_LOGIC is array ( 0 to HOLE_COUNT - 1 ) of std_logic;
	
	signal holeMinX : HOLE_ARR_UNSIGNED;
	signal holeMinY : HOLE_ARR_UNSIGNED;
	signal holeMaxX : HOLE_ARR_UNSIGNED;
	signal holeMaxY : BALL_ARR_UNSIGNED;
	signal holeOn : HOLE_ARR_LOGIC;
	
	
	signal wallRomX : integer;
	signal wallRomY : integer;
	
	signal wallR : std_logic_vector( 7 downto 0 );
	signal wallG : std_logic_vector( 7 downto 0 );
	signal wallB : std_logic_vector( 7 downto 0 );
	
	------------------------------------------------------------------------
	
	constant CUEBALL_COUNT : integer := 32;
	
    type CUEBALL_ARR_UNSIGNED is array ( 0 to CUEBALL_COUNT - 1 ) of unsigned( OBJECT_SIZE - 1 downto 0 );
    type CUEBALL_ARR_VECTOR is array ( 0 to CUEBALL_COUNT - 1 ) of std_logic_vector( 23 downto 0 );
    type CUEBALL_ARR_LOGIC is array ( 0 to CUEBALL_COUNT - 1 ) of std_logic;
	
	signal cueballMinX : CUEBALL_ARR_UNSIGNED;
	signal cueballMinY : CUEBALL_ARR_UNSIGNED;
	signal cueballMaxX : CUEBALL_ARR_UNSIGNED;
	signal cueballMaxY : CUEBALL_ARR_UNSIGNED;
	signal cueballOn : CUEBALL_ARR_LOGIC;
	
	constant addressCueballMinX : CUEBALL_ARR_UNSIGNED := (
		x"0100",
		x"0102",
		x"0104",
		x"0106",
		x"0108",
		x"010A",
		x"010C",
		x"010E",
		x"0110",
		x"0112",
		x"0114",
		x"0116",
		x"0118",
		x"011A",
		x"011C",
		x"011E",
		x"0120",
		x"0122",
		x"0124",
		x"0126",
		x"0128",
		x"012A",
		x"012C",
		x"012E",
		x"0130",
		x"0132",
		x"0134",
		x"0136",
		x"0138",
		x"013A",
		x"013C",
		x"013E"
	);
	
	constant addressCueballMinY : CUEBALL_ARR_UNSIGNED := (
		x"0101",
		x"0103",
		x"0105",
		x"0107",
		x"0109",
		x"010B",
		x"010D",
		x"010F",
		x"0111",
		x"0113",
		x"0115",
		x"0117",
		x"0119",
		x"011B",
		x"011D",
		x"011F",
		x"0121",
		x"0123",
		x"0125",
		x"0127",
		x"0129",
		x"012B",
		x"012D",
		x"012F",
		x"0131",
		x"0133",
		x"0135",
		x"0137",
		x"0139",
		x"013B",
		x"013D",
		x"013F"
	);
	
	constant cueballRgb : CUEBALL_ARR_VECTOR := (
		x"000000",
		x"FFF000",
		x"EEE000",
		x"DDD000",
		x"CCC000",
		x"BBB000",
		x"AAA000",
		x"999000",
		x"888000",
		x"777000",
		x"666000",
		x"555000",
		x"444000",
		x"333000",
		x"222000",
		x"111000",
		x"000000",
		x"000000",
		x"000000",
		x"000000",
		x"000000",
		x"000000",
		x"000000",
		x"000000",
		x"000000",
		x"000000",
		x"000000",
		x"000000",
		x"000000",
		x"000000",
		x"000000",
		x"000000"
	);
	

	-- ---------------------------------------------------------------------
	-- ---------------------------------------------------------------------
	-- ---------------------------------------------------------------------
	-- ---------------------------------------------------------------------
	-- ---------------------------------------------------------------------
	-- ---------------------------------------------------------------------
	-- ---------------------------------------------------------------------
	-- ---------------------------------------------------------------------
	-- ---------------------------------------------------------------------
	-- ---------------------------------------------------------------------

begin


	-- ---------------------------------------------------------------------
	-- ---------------------------------------------------------------------
	-- ADDED BY MAKKUS
	pixelX <= unsigned( pixel_x );
	pixelY <= unsigned( pixel_y );
	
	--varShake <= unsigned( object1x );
	varAddress <= unsigned( object2x );
	varValue <= unsigned( object2y );
	
	--
	
	--
	
	
	-- ---------------------------------------------------------------------
	-- ---------------------------------------------------------------------
	-- ---------------------------------------------------------------------



    -- draw wall and color
--    wall_on <= '1' when WALL_X_L<=pix_x and pix_x<=WALL_X_R else '0';
--    wall_rgb <= x"0000FF"; -- blue

    -- draw box and color
    -- calculate the coordinates
--    box_x_l <= unsigned(object1x);
--    box_y_t <= unsigned(object1y);
--    box_x_r <= box_x_l + BOX_SIZE_X - 1;
--    box_y_b <= box_y_t + BOX_SIZE_Y - 1;
--    box_on <= '1' when box_x_l<=pix_x and pix_x<=box_x_r and
--                      box_y_t<=pix_y and pix_y<=box_y_b else
--              '0';
    -- box rgb output
--    box_rgb <= x"00FF00"; --green

    -- draw ball and color
    -- calculate the coordinates
    
	--ball_x_l <= unsigned(object2x);
    --ball_y_t <= unsigned(object2y);
	-- MAKKUS

	--
	
	
--    ball_x_r <= ball_x_l + BALL_SIZE - 1;
--    ball_y_b <= ball_y_t + BALL_SIZE - 1;

--    square_ball_on <= '1' when ball_x_l<=pix_x and pix_x<=ball_x_r and
--                               ball_y_t<=pix_y and pix_y<=ball_y_b else
--                      '0';
    -- map current pixel location to ROM addr/col
--    rom_addr <= pix_y(2 downto 0) - ball_y_t(2 downto 0);
--    rom_col <= pix_x(2 downto 0) - ball_x_l(2 downto 0);
--    rom_bit <= BALL_ROM(to_integer(rom_addr))(to_integer(rom_col));
    -- pixel within ball
 --   ball_on <= '1' when square_ball_on='1' and rom_bit='1' else '0';
    -- ball rgb output
--    ball_rgb <= x"FF0000";   -- red

    -- display the image based on who is active
    -- note that the order is important
  --  process(video_active, wall_on, box_on, wall_rgb, box_rgb, ball_rgb, backgrnd_rgb, ball_on) is
 --   begin
--		if video_active='0' then
--			rgb <= x"000000"; --blank
--		else
--			if wall_on='1' then
--				rgb <= wall_rgb;
--			elsif ball_on='1' then
--				rgb <= ball_rgb;
--			elsif box_on='1' then
    --         rgb <= box_rgb;
    --      else
    --         rgb <= backgrnd_rgb; -- x"FFFF00"; -- yellow background
    --      end if;
    --   end if;
    --end process;
	
	-- ---------------------------------------------------------------------
	-- ---------------------------------------------------------------------
	-- ADDED BY MAKKUS
	
--	process( varAddress, varValue, ballMinX_1 ) is
--	begin
--		if varAddress = 255 then
--			ballMinX_1 <= varValue;
--		end if;
--	end process;
	
--	process( varAddress, varValue, ballMinY_1 ) is
--	begin
--		if varAddress = 254 then
--			ballMinY_1 <= varValue;
--		end if;
--	end process;
	
--	process( varAddress, varValue, ballMinX_2 ) is
--	begin
--		if varAddress = 253 then
--			ballMinX_2 <= varValue;
--		end if;
--	end process;
	
--	process( varAddress, varValue, ballMinY_2 ) is
--	begin
--		if varAddress = 252 then
--			ballMinY_2 <= varValue;
--		end if;
--	end process;
	
--	process( varAddress, varValue, ballMinX_3 ) is
--	begin
--		if varAddress = 251 then
--			ballMinX_3 <= varValue;
--		end if;
--	end process;
	
--	process( varAddress, varValue, ballMinY_3 ) is
--	begin
--		if varAddress = 250 then
--			ballMinY_3 <= varValue;
--		end if;
--	end process;

	GEN_BALL_X : for idx in 0 to BALL_COUNT - 1 generate
		process( S_AXI_ACLK ) is
		begin
			if rising_edge( S_AXI_ACLK ) then
				if varAddress = addressMinX( idx ) then
					ballMinX( idx ) <= varValue;
				end if;
			end if;
		end process;
	end generate GEN_BALL_X;

	GEN_BALL_Y : for idx in 0 to BALL_COUNT - 1 generate
		process( S_AXI_ACLK ) is
		begin
			if rising_edge( S_AXI_ACLK ) then
				if varAddress = addressMinY( idx ) then
					ballMinY( idx ) <= varValue;
				end if;
			end if;
		end process;
	end generate GEN_BALL_Y;
	
	GEN_BALL : for idx in 0 to BALL_COUNT - 1 generate
		ballMaxX( idx ) <= ballMinX( idx ) + BALL_SIZE_32 - 1;
		ballMaxY( idx ) <= ballMinY( idx ) + BALL_SIZE_32 - 1;
		ballOn( idx ) <= '1' when
			ballMinX( idx ) <= pixelX
			and pixelX <= ballMaxX( idx )
			and ballMinY( idx ) <= pixelY
			and pixelY <= ballMaxY( idx )
			and	BALL_ROM_32( to_integer( pixelY( 4 downto 0 ) - ballMinY( idx )( 4 downto 0 ) ) )( to_integer( pixelX( 4 downto 0 ) - ballMinX( idx )( 4 downto 0 ) ) ) = '1'
		else '0';
	end generate GEN_BALL;
	
	
	
	
	
	
	
	
	
	
	
	
	GEN_CUEBALL_X : for idx in 0 to CUEBALL_COUNT - 1 generate
		process( S_AXI_ACLK ) is
		begin
			if rising_edge( S_AXI_ACLK ) then
				if varAddress = addressCueballMinX( idx ) then
					cueballMinX( idx ) <= varValue;
				end if;
			end if;
		end process;
	end generate GEN_CUEBALL_X;

	GEN_CUEBALL_Y : for idx in 0 to CUEBALL_COUNT - 1 generate
		process( S_AXI_ACLK ) is
		begin
			if rising_edge( S_AXI_ACLK ) then
				if varAddress = addressCueballMinY( idx ) then
					cueballMinY( idx ) <= varValue;
				end if;
			end if;
		end process;
	end generate GEN_CUEBALL_Y;
	
	GEN_CUEBALL : for idx in 0 to CUEBALL_COUNT - 1 generate
		cueballMaxX( idx ) <= cueballMinX( idx ) + BALL_SIZE_8 - 1;
		cueballMaxY( idx ) <= cueballMinY( idx ) + BALL_SIZE_8 - 1;
		cueballOn( idx ) <= '1' when
			cueballMinX( idx ) <= pixelX
			and pixelX <= cueballMaxX( idx )
			and cueballMinY( idx ) <= pixelY
			and pixelY <= cueballMaxY( idx )
			and	BALL_ROM_8( to_integer( pixelY( 2 downto 0 ) - cueballMinY( idx )( 2 downto 0 ) ) )( to_integer( pixelX( 2 downto 0 ) - cueballMinX( idx )( 2 downto 0 ) ) ) = '1'
		else '0';
	end generate GEN_CUEBALL;
	
	
	
	
	
	
	
	
	
	
	holeMinX( 0 ) <= to_unsigned( 40 - 16 + 4, 16 );
	holeMinX( 1 ) <= to_unsigned( 640 - 16, 16 );
	holeMinX( 2 ) <= to_unsigned( ( 1240 - 16 ) - 4, 16 );
	holeMinX( 3 ) <= to_unsigned( 40 - 16 + 4, 16 );
	holeMinX( 4 ) <= to_unsigned( 640 - 16, 16 );
	holeMinX( 5 ) <= to_unsigned( ( 1240 - 16 ) - 4, 16 );
	
	holeMinY( 0 ) <= to_unsigned( 40 - 16 + 4, 16 );
	holeMinY( 1 ) <= to_unsigned( 40 - 16 + 4, 16 );
	holeMinY( 2 ) <= to_unsigned( 40 - 16 + 4, 16 );
	holeMinY( 3 ) <= to_unsigned( ( 640 - 16 ) - 4, 16 );
	holeMinY( 4 ) <= to_unsigned( ( 640 - 16 ) - 4, 16 );
	holeMinY( 5 ) <= to_unsigned( ( 640 - 16 ) - 4, 16 );
	
	GEN_HOLE : for idx in 0 to 5 generate
		holeMaxX( idx ) <= holeMinX( idx ) + BALL_SIZE_32 - 1;
		holeMaxY( idx ) <= holeMinY( idx ) + BALL_SIZE_32 - 1;
		holeOn( idx ) <= '1' when
			holeMinX( idx ) <= pixelX
			and pixelX <= holeMaxX( idx )
			and holeMinY( idx ) <= pixelY
			and pixelY <= holeMaxY( idx )
			and	BALL_ROM_32( to_integer( pixelY( 4 downto 0 ) - holeMinY( idx )( 4 downto 0 ) ) )( to_integer( pixelX( 4 downto 0 ) - holeMinX( idx )( 4 downto 0 ) ) ) = '1'
		else '0';
	end generate GEN_HOLE;
	
	
	
	
	
	
--	process( video_active, ballOn ) is
--    begin
--		ballIdx <= 0;
--		pixelIsBackground <= true;
--		for idx in 0 to BALL_COUNT - 1 loop 
--			if ballOn( idx ) = '1' then
--				ballIdx <= idx;
--				pixelIsBackground <= false;
--			end if;
--		end loop;
 --   end process;
	
	ballIdx <=
		0 when ballOn( 0 ) = '1' else
		1 when ballOn( 1 ) = '1' else
		2 when ballOn( 2 ) = '1' else
		3 when ballOn( 3 ) = '1' else
		4 when ballOn( 4 ) = '1' else
		5 when ballOn( 5 ) = '1' else
		6 when ballOn( 6 ) = '1' else
		7 when ballOn( 7 ) = '1' else
		8 when ballOn( 8 ) = '1' else
		9 when ballOn( 9 ) = '1' else
		10 when ballOn( 10 ) = '1' else
		11 when ballOn( 11 ) = '1' else
		12 when ballOn( 12 ) = '1' else
		13 when ballOn( 13 ) = '1' else
		14 when ballOn( 14 ) = '1' else
		15 when ballOn( 15 ) = '1' else
		0;
		
	cueballIdx <=
		0 when cueballOn( 0 ) = '1' else
		1 when cueballOn( 1 ) = '1' else
		2 when cueballOn( 2 ) = '1' else
		3 when cueballOn( 3 ) = '1' else
		4 when cueballOn( 4 ) = '1' else
		5 when cueballOn( 5 ) = '1' else
		6 when cueballOn( 6 ) = '1' else
		7 when cueballOn( 7 ) = '1' else
		8 when cueballOn( 8 ) = '1' else
		9 when cueballOn( 9 ) = '1' else
		10 when cueballOn( 10 ) = '1' else
		11 when cueballOn( 11 ) = '1' else
		12 when cueballOn( 12 ) = '1' else
		13 when cueballOn( 13 ) = '1' else
		14 when cueballOn( 14 ) = '1' else
		15 when cueballOn( 15 ) = '1' else
		16 when cueballOn( 16 ) = '1' else
		17 when cueballOn( 17 ) = '1' else
		18 when cueballOn( 18 ) = '1' else
		19 when cueballOn( 19 ) = '1' else
		20 when cueballOn( 20 ) = '1' else
		21 when cueballOn( 21 ) = '1' else
		22 when cueballOn( 22 ) = '1' else
		23 when cueballOn( 23 ) = '1' else
		24 when cueballOn( 24 ) = '1' else
		25 when cueballOn( 25 ) = '1' else
		26 when cueballOn( 26 ) = '1' else
		27 when cueballOn( 27 ) = '1' else
		28 when cueballOn( 28 ) = '1' else
		29 when cueballOn( 29 ) = '1' else
		30 when cueballOn( 30 ) = '1' else
		31 when cueballOn( 31 ) = '1' else
		0;
		
	pixelIsBall <=
		true when ballOn( 0 ) = '1' else
		true when ballOn( 1 ) = '1' else
		true when ballOn( 2 ) = '1' else
		true when ballOn( 3 ) = '1' else
		true when ballOn( 4 ) = '1' else
		true when ballOn( 5 ) = '1' else
		true when ballOn( 6 ) = '1' else
		true when ballOn( 7 ) = '1' else
		true when ballOn( 8 ) = '1' else
		true when ballOn( 9 ) = '1' else
		true when ballOn( 10 ) = '1' else
		true when ballOn( 11 ) = '1' else
		true when ballOn( 12 ) = '1' else
		true when ballOn( 13 ) = '1' else
		true when ballOn( 14 ) = '1' else
		true when ballOn( 15 ) = '1' else
		false;
		
	pixelIsCueball <=
		true when cueballOn( 0 ) = '1' else
		true when cueballOn( 1 ) = '1' else
		true when cueballOn( 2 ) = '1' else
		true when cueballOn( 3 ) = '1' else
		true when cueballOn( 4 ) = '1' else
		true when cueballOn( 5 ) = '1' else
		true when cueballOn( 6 ) = '1' else
		true when cueballOn( 7 ) = '1' else
		true when cueballOn( 8 ) = '1' else
		true when cueballOn( 9 ) = '1' else
		true when cueballOn( 10 ) = '1' else
		true when cueballOn( 11 ) = '1' else
		true when cueballOn( 12 ) = '1' else
		true when cueballOn( 13 ) = '1' else
		true when cueballOn( 14 ) = '1' else
		true when cueballOn( 15 ) = '1' else
		true when cueballOn( 16 ) = '1' else
		true when cueballOn( 17 ) = '1' else
		true when cueballOn( 18 ) = '1' else
		true when cueballOn( 19 ) = '1' else
		true when cueballOn( 20 ) = '1' else
		true when cueballOn( 21 ) = '1' else
		true when cueballOn( 22 ) = '1' else
		true when cueballOn( 23 ) = '1' else
		true when cueballOn( 24 ) = '1' else
		true when cueballOn( 25 ) = '1' else
		true when cueballOn( 26 ) = '1' else
		true when cueballOn( 27 ) = '1' else
		true when cueballOn( 28 ) = '1' else
		true when cueballOn( 29 ) = '1' else
		true when cueballOn( 30 ) = '1' else
		true when cueballOn( 31 ) = '1' else
		false;
		
	pixelIsHole <=
		true when holeOn( 0 ) = '1' else
		true when holeOn( 1 ) = '1' else
		true when holeOn( 2 ) = '1' else
		true when holeOn( 3 ) = '1' else
		true when holeOn( 4 ) = '1' else
		true when holeOn( 5 ) = '1' else
		false;

	
	ballR <= to_integer( unsigned( ballRgb( ballIdx )( 23 downto 16 ) ) );
	ballG <= to_integer( unsigned( ballRgb( ballIdx )( 15 downto 8 ) ) );
	ballB <= to_integer( unsigned( ballRgb( ballIdx )( 7 downto 0 ) ) );
	romX <= to_integer( pixelX( 4 downto 0 ) - ballMinX( ballIdx )( 4 downto 0 ) );
	romY <= to_integer( pixelY( 4 downto 0 ) - ballMinY( ballIdx )( 4 downto 0 ) );
	shadeR <= BALL32_COLOR( romY, romX );
	shadeG <= BALL32_COLOR( romY, romX );
	shadeB <= BALL32_COLOR( romY, romX );
	shadeA <= BALL32_ALPHA( romY, romX );
	pixR <= ( shadeR * shadeA + ( 255 - shadeA ) * ballR );
	pixG <= ( shadeG * shadeA + ( 255 - shadeA ) * ballG );
	pixB <= ( shadeB * shadeA + ( 255 - shadeA ) * ballB );
	pixVecR <= std_logic_vector( to_unsigned( pixR, 16 ) );
	pixVecG <= std_logic_vector( to_unsigned( pixG, 16 ) );
	pixVecB <= std_logic_vector( to_unsigned( pixB, 16 ) );
	
	wallRomX <= to_integer( pixelX ) mod 40;
	wallRomY <= to_integer( pixelY ) mod 40;
	pixelIsWall <= 
		pixelIsBall = false
		and
		(
			( pixelY >= 0 and pixelY < 40 and pixelX >=0 and pixelX < 1280 )
			or
			( pixelY >= 640 and pixelY < 680 and pixelX >=0 and pixelX < 1280 )
			or
			( pixelY >= 0 and pixelY < 680 and pixelX >=0 and pixelX < 40 )
			or
			( pixelY >= 0 and pixelY < 680 and pixelX >=1240 and pixelX < 1280 )
		)
	;
	wallR <= std_logic_vector( to_unsigned( WALL40_COLOR_R( wallRomY, wallRomX ), 8 ) );
	wallG <= std_logic_vector( to_unsigned( WALL40_COLOR_G( wallRomY, wallRomX ), 8 ) );
	wallB <= std_logic_vector( to_unsigned( WALL40_COLOR_B( wallRomY, wallRomX ), 8 ) );
	
	pixelIsTable <= 
		pixelIsBall = false
		and
		pixelIsWall = false
		and
		(
			( pixelY >= 0 and pixelY < 680 and pixelX >=0 and pixelX < 1280 )
		)
	;
	
	rgb( 23 downto 16 ) <=
		cueballRgb( cueballIdx )( 23 downto 16 ) when pixelIsCueball else
		pixVecR( 15 downto 8 ) when pixelIsBall else
		x"00" when pixelIsHole else
		wallR when pixelIsWall else
		x"00" when pixelIsTable else
		x"00"
	;
	
	rgb( 15 downto 8 ) <=
		cueballRgb( cueballIdx )( 15 downto 8 ) when pixelIsCueball else
		pixVecG( 15 downto 8 ) when pixelIsBall else
		x"00" when pixelIsHole else
		wallG when pixelIsWall else
		x"66" when pixelIsTable else
		x"00"
	;
	
	rgb( 7 downto 0 ) <=
		cueballRgb( cueballIdx )( 7 downto 0 ) when pixelIsCueball else
		pixVecB( 15 downto 8 ) when pixelIsBall else
		x"00" when pixelIsHole else
		wallB when pixelIsWall else
		x"00" when pixelIsTable else
		x"00"
	;
	
	-- ---------------------------------------------------------------------
	-- ---------------------------------------------------------------------
	-- ---------------------------------------------------------------------
	

end rtl;